`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Convert whatever encoding the input data type is into 2's complement
// 
//////////////////////////////////////////////////////////////////////////////////
module input_to_2comp(
    );


endmodule
